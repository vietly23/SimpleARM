module alu (input logic [31:0] a, b,
	output logic [31:0] c,
	output logic [3:0] flags)

end module
